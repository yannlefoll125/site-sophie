<?xml version="1.0" encoding="UTF-8"?>
<Batch version="2.0"><TaskList><Task type="WatermarkTextTask" enabled="True"><Text><![CDATA[Crédit photo : Christophe François]]></Text><Width WidthAuto="True">10</Width><Height HeightAuto="True">10</Height><Font FontSize="20" FontBold="True" FontItalic="False" FontUnderline="False" FontColor="#FFFFFF" FontCharset="1">Arial</Font><Transparency>100</Transparency><Operation>0</Operation><RotateAngle>0</RotateAngle><HorizontalJustification>2</HorizontalJustification><VerticalJustification>2</VerticalJustification><HorizontalOffset HorizontalOffsetUnit="0" HorizontalOffsetDir="0">0</HorizontalOffset><VerticalOffset VerticalOffsetUnit="0" VerticalOffsetDir="0">0</VerticalOffset><AddShadow>True</AddShadow></Task></TaskList></Batch>
